ARCHITECTURE studentVersion OF ahbRegulator IS
BEGIN

  -- AHB-Lite
  hRData  <=	(OTHERS => '0');
  hReady  <=	'0';	
  hResp	  <=	'0';	

  --
  
  
END ARCHITECTURE studentVersion;

